{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","jsonProperties":{"viewDetails":{}},"code":{"spec":"0x1","scope":"0x1","value":"MyView2020"},"model":"0x10","categorySelectorId":"0","displayStyleId":"0x20000000056","cameraOn":true,"origin":[706937.683679173,231313.84710078413,45.98981015563432],"extents":[60.2009048526238,28.22358408492344,30.10045242671205],"angles":{"pitch":-14.076426121769932,"roll":-73.44807892712345,"yaw":4.134357442929689},"camera":{"lens":89.99999999928959,"focusDist":30.10045242668512,"eye":[706960.3486319613,231281.55051639894,68.00794249663858]},"modelSelectorId":"0"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","code":{"spec":"0x1","scope":"0x1","value":""},"model":"0x10","categories":["0x20000000008","0x20000000041","0x20000000043","0x20000000045","0x20000000047","0x20000000049","0x2000000004b","0x2000000004d","0x2000000004f"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x20000000056","jsonProperties":{"styles":{"environment":{"sky":{"display":true,"groundColor":8228728,"zenithColor":16741686,"nadirColor":3880,"skyColor":16764303},"ground":{"display":false,"elevation":-0.01,"aboveColor":25600,"belowColor":2179941}},"hline":{"hidden":{"color":0,"ovrColor":true,"pattern":3435973836,"width":1},"transThreshold":0.3,"visible":{"color":0,"ovrColor":true,"pattern":0,"width":1}},"sceneLights":{"ambient":{"intensity":20,"type":2},"fstop":0.8570573925971985,"portrait":{"intensity":100,"intensity2":100,"type":4},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1]},"subCategoryOvr":null,"viewflags":{"renderMode":6,"noSourceLights":false,"noCameraLights":false,"noSolarLight":false,"noConstruct":true,"noTransp":false,"visEdges":false,"backgroundMap":true}}},"code":{"spec":"0xa","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","code":{"spec":"0x1","scope":"0x1","value":""},"model":"0x10","models":["0x20000000030"]}}