{"location":[706959.4849118192,231307.9950550787,57.19610878598451],"iconIndex":0,"severity":10,"id":0,"text":"信号灯放置位置不合适，请修正。"}