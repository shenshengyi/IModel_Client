{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x2000000003b","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007","categorySelectorId":"0x2000000003e","displayStyleId":"0x2000000003d","isPrivate":false,"description":"","cameraOn":true,"origin":[96645.36716324098,80510.39518881467,-1.5975356773601141],"extents":[11.090105164023587,4.876942636593589,12.839514296130522],"angles":{"pitch":-42.388753647486375,"roll":-55.4808403338392,"yaw":24.87562521004348},"camera":{"lens":46.716522041620486,"focusDist":12.839514296002688,"eye":[96640.84737038726,80498.84519401804,6.200251503494698]},"modelSelectorId":"0x2000000003c"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x2000000003e","code":{"spec":"0x8","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007","categories":["0x20000000008"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x2000000003d","jsonProperties":{"styles":{"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}},"hline":{"hidden":{"color":0,"ovrColor":true,"pattern":3435973836,"width":1},"transThreshold":0.3,"visible":{"color":0,"ovrColor":true,"pattern":0,"width":1}},"sceneLights":{"ambient":{"intensity":20,"type":2},"fstop":0.8570573925971985,"portrait":{"intensity":100,"intensity2":100,"type":4},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1]},"subCategoryOvr":null,"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true}}},"code":{"spec":"0xa","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x2000000003c","code":{"spec":"0x11","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007","models":["0x20000000030"]}}