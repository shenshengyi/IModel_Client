{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","jsonProperties":{"viewDetails":{}},"code":{"spec":"0x1","scope":"0x1","value":"MyView2020"},"model":"0x10","categorySelectorId":"0","displayStyleId":"0x2000000003d","cameraOn":true,"origin":[96644.88442283828,80510.42728846685,-48.283022056270255],"extents":[216.6393055920489,101.56554411254051,3.3711281822616],"angles":{"roll":-90},"camera":{"lens":90,"focusDist":108.31965279602447,"eye":[96753.2040756343,80398.73650748856,2.49975]},"modelSelectorId":"0"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","code":{"spec":"0x1","scope":"0x1","value":""},"model":"0x10","categories":["0x20000000008","0x40000000002","0x40000000006","0x4000000000a","0x4000000000e","0x40000000012","0x40000000016","0x4000000001a","0x4000000001e","0x40000000022","0x40000000026","0x4000000002a","0x4000000002e","0x40000000032","0x40000000036","0x4000000003a","0x4000000003e","0x40000000042","0x40000000046","0x4000000004a","0x4000000004e","0x40000000052","0x40000000056","0x4000000005a","0x4000000005e","0x40000000062","0x40000000066","0x4000000006a","0x4000000006e","0x40000000072","0x40000000076","0x4000000007a","0x4000000007e","0x40000000082","0x40000000086","0x4000000008a","0x4000000008e","0x40000000092","0x40000000096","0x4000000009a","0x4000000009e","0x400000000a2","0x400000000a6","0x400000000aa","0x400000000ae","0x400000000b2","0x400000000b6","0x400000000ba","0x400000000be","0x400000000c2","0x400000000c6","0x400000000ca","0x400000000ce","0x400000000d2","0x400000000d6","0x400000000da","0x400000000de","0x400000000e2","0x400000000f2","0x400000000f6","0x400000000fa","0x40000000101","0x40000000105","0x40000000109","0x4000000010d","0x40000000111","0x40000000113","0x40000000118","0x4000000011a","0x4000000011f","0x40000000121","0x40000000126","0x40000000128","0x4000000012d","0x4000000012f","0x40000000134","0x40000000136","0x4000000013b","0x4000000013f","0x40000000143","0x40000000145","0x4000000014a","0x4000000014c","0x40000000151","0x40000000153","0x40000000158","0x4000000015a","0x4000000015f","0x40000000161","0x40000000166","0x40000000168","0x4000000016d","0x40000000171","0x40000000175","0x40000000179","0x4000000017d","0x40000000181","0x40000000185","0x40000000189","0x4000000018d","0x40000000191","0x40000000195","0x40000000199","0x4000000019d","0x400000001a1","0x400000001a5","0x400000001a9","0x400000001ad","0x400000001b1","0x400000001b5","0x400000001b9","0x400000001bd","0x400000001c1","0x400000001c5","0x400000001c9","0x400000001cd","0x400000001d1","0x400000001d5","0x400000001d9","0x400000001dd","0x400000001e1","0x400000001ed","0x400000001f5","0x40000000201","0x40000000205","0x40000000211","0x40000000215","0x4000000021d","0x40000000221","0x4000000022d","0x40000000231","0x40000000235","0x40000000239","0x40000000245","0x40000000275","0x40000000279","0x40000000285","0x4000000028d","0x40000000299","0x4000000029d","0x400000002a1","0x400000002b1","0x400000002c1","0x400000002c5"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x2000000003d","jsonProperties":{"styles":{"environment":{"sky":{"display":true,"groundColor":8228728,"zenithColor":16741686,"nadirColor":3880,"skyColor":16764303},"ground":{"display":false,"elevation":-0.01,"aboveColor":25600,"belowColor":2179941}},"hline":{"hidden":{"color":0,"ovrColor":true,"pattern":3435973836,"width":1},"transThreshold":0.3,"visible":{"color":0,"ovrColor":true,"pattern":0,"width":1}},"sceneLights":{"ambient":{"intensity":20,"type":2},"fstop":0.8570573925971985,"portrait":{"intensity":100,"intensity2":100,"type":4},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1]},"subCategoryOvr":null,"viewflags":{"renderMode":6,"noSourceLights":false,"noCameraLights":false,"noSolarLight":false,"noConstruct":true,"noTransp":false,"visEdges":false,"backgroundMap":true}}},"code":{"spec":"0xa","scope":"0x20000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x20000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","code":{"spec":"0x1","scope":"0x1","value":""},"model":"0x10","models":["0x400000002c4","0x400000002c0","0x400000002bc","0x400000002b8","0x400000002b4","0x400000002b0","0x400000002ac","0x400000002a8","0x400000002a4","0x400000002a0","0x4000000029c","0x40000000298","0x40000000294","0x40000000290","0x4000000028c","0x40000000288","0x40000000284","0x40000000280","0x4000000027c","0x40000000278","0x40000000274","0x40000000270","0x4000000026c","0x40000000268","0x40000000264","0x40000000260","0x4000000025c","0x40000000258","0x40000000254","0x40000000250","0x4000000024c","0x40000000248","0x40000000244","0x40000000240","0x4000000023c","0x40000000238","0x40000000234","0x40000000230","0x4000000022c","0x40000000228","0x40000000224","0x40000000220","0x4000000021c","0x40000000218","0x40000000214","0x40000000210","0x4000000020c","0x40000000208","0x40000000204","0x40000000200","0x400000001fc","0x400000001f8","0x400000001f4","0x400000001f0","0x400000001ec","0x400000001e8","0x400000001e4","0x20000000030"]}}